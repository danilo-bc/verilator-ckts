module and_custom(input A,
                  input B,
                  
                  output S);

    assign S = A&B;
endmodule
    
